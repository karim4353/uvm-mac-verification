`timescale 1ns/1ps
module random_stress_test;
    initial begin
        $display("Random stress test placeholder - run under Questa/Xcelium for UVM sequences");
        #10 $finish;
    end
endmodule
