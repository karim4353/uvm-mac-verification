package uvm_mac_pkg;
    import uvm_pkg::*;
    // covergroup placeholders
    covergroup cg_packet_size;
        option.per_instance = 1;
        size: coverpoint int'(0);
    endgroup
endpackage
